library verilog;
use verilog.vl_types.all;
entity ins_decoder is
    port(
        instruction     : in     vl_logic_vector(42 downto 0);
        dec_src_dat_ram_addr_en_b: out    vl_logic;
        dec_src_dat_ram_addr: out    vl_logic_vector(16 downto 0);
        dec_src_imm_dat_sel: out    vl_logic;
        dec_src_imm_dat : out    vl_logic_vector(15 downto 0);
        dec_src_indir_addr_sel: out    vl_logic;
        dec_src_r0_r_sel: out    vl_logic;
        dec_src_r1_r_sel: out    vl_logic;
        dec_src_r2_r_sel: out    vl_logic;
        dec_src_r3_r_sel: out    vl_logic;
        dec_src_r4_r_sel: out    vl_logic;
        dec_src_r5_r_sel: out    vl_logic;
        dec_src_r6_r_sel: out    vl_logic;
        dec_src_r7_r_sel: out    vl_logic;
        dec_src_sprf0_r_sel: out    vl_logic;
        dec_src_sprf1_r_sel: out    vl_logic;
        dec_src_r0_t_sel: out    vl_logic;
        dec_src_r1_t_sel: out    vl_logic;
        dec_src_r2_t_sel: out    vl_logic;
        dec_src_r3_t_sel: out    vl_logic;
        dec_src_r4_t_sel: out    vl_logic;
        dec_src_r5_t_sel: out    vl_logic;
        dec_src_r6_t_sel: out    vl_logic;
        dec_src_r7_t_sel: out    vl_logic;
        dec_src_rmod_t_sel: out    vl_logic;
        dec_dst_dat_ram_addr_en_b: out    vl_logic;
        dec_dst_dat_ram_rw: out    vl_logic;
        dec_dst_dat_ram_addr: out    vl_logic_vector(16 downto 0);
        dec_dst_indir_addr_sel: out    vl_logic;
        dec_dst_r0_r_sel: out    vl_logic;
        dec_dst_r1_r_sel: out    vl_logic;
        dec_dst_r2_r_sel: out    vl_logic;
        dec_dst_r3_r_sel: out    vl_logic;
        dec_dst_r4_r_sel: out    vl_logic;
        dec_dst_r5_r_sel: out    vl_logic;
        dec_dst_r6_r_sel: out    vl_logic;
        dec_dst_r7_r_sel: out    vl_logic;
        dec_dst_sprf0_r_sel: out    vl_logic;
        dec_dst_sprf1_r_sel: out    vl_logic;
        dec_dst_r0_t_sel: out    vl_logic;
        dec_dst_r1_t_sel: out    vl_logic;
        dec_dst_r2_t_sel: out    vl_logic;
        dec_dst_r3_t_sel: out    vl_logic;
        dec_dst_r4_t_sel: out    vl_logic;
        dec_dst_r5_t_sel: out    vl_logic;
        dec_dst_r6_t_sel: out    vl_logic;
        dec_dst_r7_t_sel: out    vl_logic;
        dec_dst_rmod_t_sel: out    vl_logic;
        dec_dst_jmp_addr_sel: out    vl_logic;
        dec_dst_jmp_addr: out    vl_logic_vector(18 downto 0);
        dec_opr_typ_sel : out    vl_logic_vector(4 downto 0);
        dec_opr_div_mod_sel: out    vl_logic;
        dec_alu_o_sel   : out    vl_logic;
        dec_alu_t_sel   : out    vl_logic;
        dec_alu_typ_sel : out    vl_logic_vector(3 downto 0);
        dec_prng_t_sel  : out    vl_logic;
        dec_prng_typ_sel: out    vl_logic_vector(1 downto 0);
        dec_sprf_r0_typ_sel: out    vl_logic_vector(1 downto 0);
        dec_sprf_r1_typ_sel: out    vl_logic_vector(1 downto 0);
        dec_delay_src_dst_sel: out    vl_logic;
        dec_delay_src_dst: out    vl_logic_vector(7 downto 0)
    );
end ins_decoder;
