library verilog;
use verilog.vl_types.all;
entity MUL_32bit_tb is
    generic(
        n               : integer := 32
    );
end MUL_32bit_tb;
