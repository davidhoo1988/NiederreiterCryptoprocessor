library verilog;
use verilog.vl_types.all;
entity gopf_mul_tb is
end gopf_mul_tb;
