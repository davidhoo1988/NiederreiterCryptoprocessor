library verilog;
use verilog.vl_types.all;
entity split_tb is
end split_tb;
